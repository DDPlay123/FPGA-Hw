// NIOS_LED_Qsys.v

// Generated using ACDS version 18.1 625

`timescale 1 ps / 1 ps
module NIOS_LED_Qsys (
		input  wire       clk_clk,                        //                     clk.clk
		output wire [7:0] led_external_connection_export, // led_external_connection.export
		input  wire       reset_reset_n,                  //                   reset.reset_n
		input  wire       sw_external_connection_export   //  sw_external_connection.export
	);

	wire         pll_outclk0_clk;                                             // pll:outclk_0 -> [NIOS_CPU:clk, irq_mapper:clk, irq_synchronizer:sender_clk, irq_synchronizer_001:sender_clk, jtag_uart:clk, mm_interconnect_0:pll_outclk0_clk, mm_interconnect_1:pll_outclk0_clk, onchip_memory:clk, rst_controller_001:clk]
	wire         pll_outclk1_clk;                                             // pll:outclk_1 -> [LED:clk, SW:clk, irq_synchronizer:receiver_clk, irq_synchronizer_001:receiver_clk, mm_clock_crossing_bridge:m0_clk, mm_clock_crossing_bridge:s0_clk, mm_interconnect_0:pll_outclk1_clk, mm_interconnect_1:pll_outclk1_clk, rst_controller:clk, rst_controller_002:clk, sysid:clock, timer_10ms:clk, timer_1ms:clk]
	wire  [31:0] nios_cpu_data_master_readdata;                               // mm_interconnect_0:NIOS_CPU_data_master_readdata -> NIOS_CPU:d_readdata
	wire         nios_cpu_data_master_waitrequest;                            // mm_interconnect_0:NIOS_CPU_data_master_waitrequest -> NIOS_CPU:d_waitrequest
	wire         nios_cpu_data_master_debugaccess;                            // NIOS_CPU:debug_mem_slave_debugaccess_to_roms -> mm_interconnect_0:NIOS_CPU_data_master_debugaccess
	wire  [24:0] nios_cpu_data_master_address;                                // NIOS_CPU:d_address -> mm_interconnect_0:NIOS_CPU_data_master_address
	wire   [3:0] nios_cpu_data_master_byteenable;                             // NIOS_CPU:d_byteenable -> mm_interconnect_0:NIOS_CPU_data_master_byteenable
	wire         nios_cpu_data_master_read;                                   // NIOS_CPU:d_read -> mm_interconnect_0:NIOS_CPU_data_master_read
	wire         nios_cpu_data_master_write;                                  // NIOS_CPU:d_write -> mm_interconnect_0:NIOS_CPU_data_master_write
	wire  [31:0] nios_cpu_data_master_writedata;                              // NIOS_CPU:d_writedata -> mm_interconnect_0:NIOS_CPU_data_master_writedata
	wire  [31:0] nios_cpu_instruction_master_readdata;                        // mm_interconnect_0:NIOS_CPU_instruction_master_readdata -> NIOS_CPU:i_readdata
	wire         nios_cpu_instruction_master_waitrequest;                     // mm_interconnect_0:NIOS_CPU_instruction_master_waitrequest -> NIOS_CPU:i_waitrequest
	wire  [24:0] nios_cpu_instruction_master_address;                         // NIOS_CPU:i_address -> mm_interconnect_0:NIOS_CPU_instruction_master_address
	wire         nios_cpu_instruction_master_read;                            // NIOS_CPU:i_read -> mm_interconnect_0:NIOS_CPU_instruction_master_read
	wire  [31:0] mm_interconnect_0_nios_cpu_debug_mem_slave_readdata;         // NIOS_CPU:debug_mem_slave_readdata -> mm_interconnect_0:NIOS_CPU_debug_mem_slave_readdata
	wire         mm_interconnect_0_nios_cpu_debug_mem_slave_waitrequest;      // NIOS_CPU:debug_mem_slave_waitrequest -> mm_interconnect_0:NIOS_CPU_debug_mem_slave_waitrequest
	wire         mm_interconnect_0_nios_cpu_debug_mem_slave_debugaccess;      // mm_interconnect_0:NIOS_CPU_debug_mem_slave_debugaccess -> NIOS_CPU:debug_mem_slave_debugaccess
	wire   [8:0] mm_interconnect_0_nios_cpu_debug_mem_slave_address;          // mm_interconnect_0:NIOS_CPU_debug_mem_slave_address -> NIOS_CPU:debug_mem_slave_address
	wire         mm_interconnect_0_nios_cpu_debug_mem_slave_read;             // mm_interconnect_0:NIOS_CPU_debug_mem_slave_read -> NIOS_CPU:debug_mem_slave_read
	wire   [3:0] mm_interconnect_0_nios_cpu_debug_mem_slave_byteenable;       // mm_interconnect_0:NIOS_CPU_debug_mem_slave_byteenable -> NIOS_CPU:debug_mem_slave_byteenable
	wire         mm_interconnect_0_nios_cpu_debug_mem_slave_write;            // mm_interconnect_0:NIOS_CPU_debug_mem_slave_write -> NIOS_CPU:debug_mem_slave_write
	wire  [31:0] mm_interconnect_0_nios_cpu_debug_mem_slave_writedata;        // mm_interconnect_0:NIOS_CPU_debug_mem_slave_writedata -> NIOS_CPU:debug_mem_slave_writedata
	wire  [31:0] mm_interconnect_0_mm_clock_crossing_bridge_s0_readdata;      // mm_clock_crossing_bridge:s0_readdata -> mm_interconnect_0:mm_clock_crossing_bridge_s0_readdata
	wire         mm_interconnect_0_mm_clock_crossing_bridge_s0_waitrequest;   // mm_clock_crossing_bridge:s0_waitrequest -> mm_interconnect_0:mm_clock_crossing_bridge_s0_waitrequest
	wire         mm_interconnect_0_mm_clock_crossing_bridge_s0_debugaccess;   // mm_interconnect_0:mm_clock_crossing_bridge_s0_debugaccess -> mm_clock_crossing_bridge:s0_debugaccess
	wire   [9:0] mm_interconnect_0_mm_clock_crossing_bridge_s0_address;       // mm_interconnect_0:mm_clock_crossing_bridge_s0_address -> mm_clock_crossing_bridge:s0_address
	wire         mm_interconnect_0_mm_clock_crossing_bridge_s0_read;          // mm_interconnect_0:mm_clock_crossing_bridge_s0_read -> mm_clock_crossing_bridge:s0_read
	wire   [3:0] mm_interconnect_0_mm_clock_crossing_bridge_s0_byteenable;    // mm_interconnect_0:mm_clock_crossing_bridge_s0_byteenable -> mm_clock_crossing_bridge:s0_byteenable
	wire         mm_interconnect_0_mm_clock_crossing_bridge_s0_readdatavalid; // mm_clock_crossing_bridge:s0_readdatavalid -> mm_interconnect_0:mm_clock_crossing_bridge_s0_readdatavalid
	wire         mm_interconnect_0_mm_clock_crossing_bridge_s0_write;         // mm_interconnect_0:mm_clock_crossing_bridge_s0_write -> mm_clock_crossing_bridge:s0_write
	wire  [31:0] mm_interconnect_0_mm_clock_crossing_bridge_s0_writedata;     // mm_interconnect_0:mm_clock_crossing_bridge_s0_writedata -> mm_clock_crossing_bridge:s0_writedata
	wire   [0:0] mm_interconnect_0_mm_clock_crossing_bridge_s0_burstcount;    // mm_interconnect_0:mm_clock_crossing_bridge_s0_burstcount -> mm_clock_crossing_bridge:s0_burstcount
	wire         mm_interconnect_0_onchip_memory_s1_chipselect;               // mm_interconnect_0:onchip_memory_s1_chipselect -> onchip_memory:chipselect
	wire  [31:0] mm_interconnect_0_onchip_memory_s1_readdata;                 // onchip_memory:readdata -> mm_interconnect_0:onchip_memory_s1_readdata
	wire  [12:0] mm_interconnect_0_onchip_memory_s1_address;                  // mm_interconnect_0:onchip_memory_s1_address -> onchip_memory:address
	wire   [3:0] mm_interconnect_0_onchip_memory_s1_byteenable;               // mm_interconnect_0:onchip_memory_s1_byteenable -> onchip_memory:byteenable
	wire         mm_interconnect_0_onchip_memory_s1_write;                    // mm_interconnect_0:onchip_memory_s1_write -> onchip_memory:write
	wire  [31:0] mm_interconnect_0_onchip_memory_s1_writedata;                // mm_interconnect_0:onchip_memory_s1_writedata -> onchip_memory:writedata
	wire         mm_interconnect_0_onchip_memory_s1_clken;                    // mm_interconnect_0:onchip_memory_s1_clken -> onchip_memory:clken
	wire         mm_clock_crossing_bridge_m0_waitrequest;                     // mm_interconnect_1:mm_clock_crossing_bridge_m0_waitrequest -> mm_clock_crossing_bridge:m0_waitrequest
	wire  [31:0] mm_clock_crossing_bridge_m0_readdata;                        // mm_interconnect_1:mm_clock_crossing_bridge_m0_readdata -> mm_clock_crossing_bridge:m0_readdata
	wire         mm_clock_crossing_bridge_m0_debugaccess;                     // mm_clock_crossing_bridge:m0_debugaccess -> mm_interconnect_1:mm_clock_crossing_bridge_m0_debugaccess
	wire   [9:0] mm_clock_crossing_bridge_m0_address;                         // mm_clock_crossing_bridge:m0_address -> mm_interconnect_1:mm_clock_crossing_bridge_m0_address
	wire         mm_clock_crossing_bridge_m0_read;                            // mm_clock_crossing_bridge:m0_read -> mm_interconnect_1:mm_clock_crossing_bridge_m0_read
	wire   [3:0] mm_clock_crossing_bridge_m0_byteenable;                      // mm_clock_crossing_bridge:m0_byteenable -> mm_interconnect_1:mm_clock_crossing_bridge_m0_byteenable
	wire         mm_clock_crossing_bridge_m0_readdatavalid;                   // mm_interconnect_1:mm_clock_crossing_bridge_m0_readdatavalid -> mm_clock_crossing_bridge:m0_readdatavalid
	wire  [31:0] mm_clock_crossing_bridge_m0_writedata;                       // mm_clock_crossing_bridge:m0_writedata -> mm_interconnect_1:mm_clock_crossing_bridge_m0_writedata
	wire         mm_clock_crossing_bridge_m0_write;                           // mm_clock_crossing_bridge:m0_write -> mm_interconnect_1:mm_clock_crossing_bridge_m0_write
	wire   [0:0] mm_clock_crossing_bridge_m0_burstcount;                      // mm_clock_crossing_bridge:m0_burstcount -> mm_interconnect_1:mm_clock_crossing_bridge_m0_burstcount
	wire         mm_interconnect_1_jtag_uart_avalon_jtag_slave_chipselect;    // mm_interconnect_1:jtag_uart_avalon_jtag_slave_chipselect -> jtag_uart:av_chipselect
	wire  [31:0] mm_interconnect_1_jtag_uart_avalon_jtag_slave_readdata;      // jtag_uart:av_readdata -> mm_interconnect_1:jtag_uart_avalon_jtag_slave_readdata
	wire         mm_interconnect_1_jtag_uart_avalon_jtag_slave_waitrequest;   // jtag_uart:av_waitrequest -> mm_interconnect_1:jtag_uart_avalon_jtag_slave_waitrequest
	wire   [0:0] mm_interconnect_1_jtag_uart_avalon_jtag_slave_address;       // mm_interconnect_1:jtag_uart_avalon_jtag_slave_address -> jtag_uart:av_address
	wire         mm_interconnect_1_jtag_uart_avalon_jtag_slave_read;          // mm_interconnect_1:jtag_uart_avalon_jtag_slave_read -> jtag_uart:av_read_n
	wire         mm_interconnect_1_jtag_uart_avalon_jtag_slave_write;         // mm_interconnect_1:jtag_uart_avalon_jtag_slave_write -> jtag_uart:av_write_n
	wire  [31:0] mm_interconnect_1_jtag_uart_avalon_jtag_slave_writedata;     // mm_interconnect_1:jtag_uart_avalon_jtag_slave_writedata -> jtag_uart:av_writedata
	wire  [31:0] mm_interconnect_1_sysid_control_slave_readdata;              // sysid:readdata -> mm_interconnect_1:sysid_control_slave_readdata
	wire   [0:0] mm_interconnect_1_sysid_control_slave_address;               // mm_interconnect_1:sysid_control_slave_address -> sysid:address
	wire  [31:0] mm_interconnect_1_sw_s1_readdata;                            // SW:readdata -> mm_interconnect_1:SW_s1_readdata
	wire   [1:0] mm_interconnect_1_sw_s1_address;                             // mm_interconnect_1:SW_s1_address -> SW:address
	wire         mm_interconnect_1_led_s1_chipselect;                         // mm_interconnect_1:LED_s1_chipselect -> LED:chipselect
	wire  [31:0] mm_interconnect_1_led_s1_readdata;                           // LED:readdata -> mm_interconnect_1:LED_s1_readdata
	wire   [1:0] mm_interconnect_1_led_s1_address;                            // mm_interconnect_1:LED_s1_address -> LED:address
	wire         mm_interconnect_1_led_s1_write;                              // mm_interconnect_1:LED_s1_write -> LED:write_n
	wire  [31:0] mm_interconnect_1_led_s1_writedata;                          // mm_interconnect_1:LED_s1_writedata -> LED:writedata
	wire         mm_interconnect_1_timer_10ms_s1_chipselect;                  // mm_interconnect_1:timer_10ms_s1_chipselect -> timer_10ms:chipselect
	wire  [15:0] mm_interconnect_1_timer_10ms_s1_readdata;                    // timer_10ms:readdata -> mm_interconnect_1:timer_10ms_s1_readdata
	wire   [2:0] mm_interconnect_1_timer_10ms_s1_address;                     // mm_interconnect_1:timer_10ms_s1_address -> timer_10ms:address
	wire         mm_interconnect_1_timer_10ms_s1_write;                       // mm_interconnect_1:timer_10ms_s1_write -> timer_10ms:write_n
	wire  [15:0] mm_interconnect_1_timer_10ms_s1_writedata;                   // mm_interconnect_1:timer_10ms_s1_writedata -> timer_10ms:writedata
	wire         mm_interconnect_1_timer_1ms_s1_chipselect;                   // mm_interconnect_1:timer_1ms_s1_chipselect -> timer_1ms:chipselect
	wire  [15:0] mm_interconnect_1_timer_1ms_s1_readdata;                     // timer_1ms:readdata -> mm_interconnect_1:timer_1ms_s1_readdata
	wire   [2:0] mm_interconnect_1_timer_1ms_s1_address;                      // mm_interconnect_1:timer_1ms_s1_address -> timer_1ms:address
	wire         mm_interconnect_1_timer_1ms_s1_write;                        // mm_interconnect_1:timer_1ms_s1_write -> timer_1ms:write_n
	wire  [15:0] mm_interconnect_1_timer_1ms_s1_writedata;                    // mm_interconnect_1:timer_1ms_s1_writedata -> timer_1ms:writedata
	wire         irq_mapper_receiver2_irq;                                    // jtag_uart:av_irq -> irq_mapper:receiver2_irq
	wire  [31:0] nios_cpu_irq_irq;                                            // irq_mapper:sender_irq -> NIOS_CPU:irq
	wire         irq_mapper_receiver0_irq;                                    // irq_synchronizer:sender_irq -> irq_mapper:receiver0_irq
	wire   [0:0] irq_synchronizer_receiver_irq;                               // timer_1ms:irq -> irq_synchronizer:receiver_irq
	wire         irq_mapper_receiver1_irq;                                    // irq_synchronizer_001:sender_irq -> irq_mapper:receiver1_irq
	wire   [0:0] irq_synchronizer_001_receiver_irq;                           // timer_10ms:irq -> irq_synchronizer_001:receiver_irq
	wire         rst_controller_reset_out_reset;                              // rst_controller:reset_out -> [LED:reset_n, mm_interconnect_1:LED_reset_reset_bridge_in_reset_reset]
	wire         nios_cpu_debug_reset_request_reset;                          // NIOS_CPU:debug_reset_request -> [rst_controller:reset_in0, rst_controller_001:reset_in1, rst_controller_002:reset_in1]
	wire         rst_controller_001_reset_out_reset;                          // rst_controller_001:reset_out -> [NIOS_CPU:reset_n, irq_mapper:reset, irq_synchronizer:sender_reset, irq_synchronizer_001:sender_reset, jtag_uart:rst_n, mm_interconnect_0:NIOS_CPU_reset_reset_bridge_in_reset_reset, mm_interconnect_1:jtag_uart_reset_reset_bridge_in_reset_reset, onchip_memory:reset, rst_translator:in_reset]
	wire         rst_controller_001_reset_out_reset_req;                      // rst_controller_001:reset_req -> [NIOS_CPU:reset_req, onchip_memory:reset_req, rst_translator:reset_req_in]
	wire         rst_controller_002_reset_out_reset;                          // rst_controller_002:reset_out -> [SW:reset_n, irq_synchronizer:receiver_reset, irq_synchronizer_001:receiver_reset, mm_clock_crossing_bridge:m0_reset, mm_clock_crossing_bridge:s0_reset, mm_interconnect_0:mm_clock_crossing_bridge_s0_reset_reset_bridge_in_reset_reset, mm_interconnect_1:mm_clock_crossing_bridge_m0_reset_reset_bridge_in_reset_reset, sysid:reset_n, timer_10ms:reset_n, timer_1ms:reset_n]

	NIOS_LED_Qsys_LED led (
		.clk        (pll_outclk1_clk),                     //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),     //               reset.reset_n
		.address    (mm_interconnect_1_led_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_1_led_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_1_led_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_1_led_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_1_led_s1_readdata),   //                    .readdata
		.out_port   (led_external_connection_export)       // external_connection.export
	);

	NIOS_LED_Qsys_NIOS_CPU nios_cpu (
		.clk                                 (pll_outclk0_clk),                                        //                       clk.clk
		.reset_n                             (~rst_controller_001_reset_out_reset),                    //                     reset.reset_n
		.reset_req                           (rst_controller_001_reset_out_reset_req),                 //                          .reset_req
		.d_address                           (nios_cpu_data_master_address),                           //               data_master.address
		.d_byteenable                        (nios_cpu_data_master_byteenable),                        //                          .byteenable
		.d_read                              (nios_cpu_data_master_read),                              //                          .read
		.d_readdata                          (nios_cpu_data_master_readdata),                          //                          .readdata
		.d_waitrequest                       (nios_cpu_data_master_waitrequest),                       //                          .waitrequest
		.d_write                             (nios_cpu_data_master_write),                             //                          .write
		.d_writedata                         (nios_cpu_data_master_writedata),                         //                          .writedata
		.debug_mem_slave_debugaccess_to_roms (nios_cpu_data_master_debugaccess),                       //                          .debugaccess
		.i_address                           (nios_cpu_instruction_master_address),                    //        instruction_master.address
		.i_read                              (nios_cpu_instruction_master_read),                       //                          .read
		.i_readdata                          (nios_cpu_instruction_master_readdata),                   //                          .readdata
		.i_waitrequest                       (nios_cpu_instruction_master_waitrequest),                //                          .waitrequest
		.irq                                 (nios_cpu_irq_irq),                                       //                       irq.irq
		.debug_reset_request                 (nios_cpu_debug_reset_request_reset),                     //       debug_reset_request.reset
		.debug_mem_slave_address             (mm_interconnect_0_nios_cpu_debug_mem_slave_address),     //           debug_mem_slave.address
		.debug_mem_slave_byteenable          (mm_interconnect_0_nios_cpu_debug_mem_slave_byteenable),  //                          .byteenable
		.debug_mem_slave_debugaccess         (mm_interconnect_0_nios_cpu_debug_mem_slave_debugaccess), //                          .debugaccess
		.debug_mem_slave_read                (mm_interconnect_0_nios_cpu_debug_mem_slave_read),        //                          .read
		.debug_mem_slave_readdata            (mm_interconnect_0_nios_cpu_debug_mem_slave_readdata),    //                          .readdata
		.debug_mem_slave_waitrequest         (mm_interconnect_0_nios_cpu_debug_mem_slave_waitrequest), //                          .waitrequest
		.debug_mem_slave_write               (mm_interconnect_0_nios_cpu_debug_mem_slave_write),       //                          .write
		.debug_mem_slave_writedata           (mm_interconnect_0_nios_cpu_debug_mem_slave_writedata),   //                          .writedata
		.dummy_ci_port                       ()                                                        // custom_instruction_master.readra
	);

	NIOS_LED_Qsys_SW sw (
		.clk      (pll_outclk1_clk),                     //                 clk.clk
		.reset_n  (~rst_controller_002_reset_out_reset), //               reset.reset_n
		.address  (mm_interconnect_1_sw_s1_address),     //                  s1.address
		.readdata (mm_interconnect_1_sw_s1_readdata),    //                    .readdata
		.in_port  (sw_external_connection_export)        // external_connection.export
	);

	NIOS_LED_Qsys_jtag_uart jtag_uart (
		.clk            (pll_outclk0_clk),                                           //               clk.clk
		.rst_n          (~rst_controller_001_reset_out_reset),                       //             reset.reset_n
		.av_chipselect  (mm_interconnect_1_jtag_uart_avalon_jtag_slave_chipselect),  // avalon_jtag_slave.chipselect
		.av_address     (mm_interconnect_1_jtag_uart_avalon_jtag_slave_address),     //                  .address
		.av_read_n      (~mm_interconnect_1_jtag_uart_avalon_jtag_slave_read),       //                  .read_n
		.av_readdata    (mm_interconnect_1_jtag_uart_avalon_jtag_slave_readdata),    //                  .readdata
		.av_write_n     (~mm_interconnect_1_jtag_uart_avalon_jtag_slave_write),      //                  .write_n
		.av_writedata   (mm_interconnect_1_jtag_uart_avalon_jtag_slave_writedata),   //                  .writedata
		.av_waitrequest (mm_interconnect_1_jtag_uart_avalon_jtag_slave_waitrequest), //                  .waitrequest
		.av_irq         (irq_mapper_receiver2_irq)                                   //               irq.irq
	);

	altera_avalon_mm_clock_crossing_bridge #(
		.DATA_WIDTH          (32),
		.SYMBOL_WIDTH        (8),
		.HDL_ADDR_WIDTH      (10),
		.BURSTCOUNT_WIDTH    (1),
		.COMMAND_FIFO_DEPTH  (32),
		.RESPONSE_FIFO_DEPTH (8),
		.MASTER_SYNC_DEPTH   (3),
		.SLAVE_SYNC_DEPTH    (3)
	) mm_clock_crossing_bridge (
		.m0_clk           (pll_outclk1_clk),                                             //   m0_clk.clk
		.m0_reset         (rst_controller_002_reset_out_reset),                          // m0_reset.reset
		.s0_clk           (pll_outclk1_clk),                                             //   s0_clk.clk
		.s0_reset         (rst_controller_002_reset_out_reset),                          // s0_reset.reset
		.s0_waitrequest   (mm_interconnect_0_mm_clock_crossing_bridge_s0_waitrequest),   //       s0.waitrequest
		.s0_readdata      (mm_interconnect_0_mm_clock_crossing_bridge_s0_readdata),      //         .readdata
		.s0_readdatavalid (mm_interconnect_0_mm_clock_crossing_bridge_s0_readdatavalid), //         .readdatavalid
		.s0_burstcount    (mm_interconnect_0_mm_clock_crossing_bridge_s0_burstcount),    //         .burstcount
		.s0_writedata     (mm_interconnect_0_mm_clock_crossing_bridge_s0_writedata),     //         .writedata
		.s0_address       (mm_interconnect_0_mm_clock_crossing_bridge_s0_address),       //         .address
		.s0_write         (mm_interconnect_0_mm_clock_crossing_bridge_s0_write),         //         .write
		.s0_read          (mm_interconnect_0_mm_clock_crossing_bridge_s0_read),          //         .read
		.s0_byteenable    (mm_interconnect_0_mm_clock_crossing_bridge_s0_byteenable),    //         .byteenable
		.s0_debugaccess   (mm_interconnect_0_mm_clock_crossing_bridge_s0_debugaccess),   //         .debugaccess
		.m0_waitrequest   (mm_clock_crossing_bridge_m0_waitrequest),                     //       m0.waitrequest
		.m0_readdata      (mm_clock_crossing_bridge_m0_readdata),                        //         .readdata
		.m0_readdatavalid (mm_clock_crossing_bridge_m0_readdatavalid),                   //         .readdatavalid
		.m0_burstcount    (mm_clock_crossing_bridge_m0_burstcount),                      //         .burstcount
		.m0_writedata     (mm_clock_crossing_bridge_m0_writedata),                       //         .writedata
		.m0_address       (mm_clock_crossing_bridge_m0_address),                         //         .address
		.m0_write         (mm_clock_crossing_bridge_m0_write),                           //         .write
		.m0_read          (mm_clock_crossing_bridge_m0_read),                            //         .read
		.m0_byteenable    (mm_clock_crossing_bridge_m0_byteenable),                      //         .byteenable
		.m0_debugaccess   (mm_clock_crossing_bridge_m0_debugaccess)                      //         .debugaccess
	);

	NIOS_LED_Qsys_onchip_memory onchip_memory (
		.clk        (pll_outclk0_clk),                               //   clk1.clk
		.address    (mm_interconnect_0_onchip_memory_s1_address),    //     s1.address
		.clken      (mm_interconnect_0_onchip_memory_s1_clken),      //       .clken
		.chipselect (mm_interconnect_0_onchip_memory_s1_chipselect), //       .chipselect
		.write      (mm_interconnect_0_onchip_memory_s1_write),      //       .write
		.readdata   (mm_interconnect_0_onchip_memory_s1_readdata),   //       .readdata
		.writedata  (mm_interconnect_0_onchip_memory_s1_writedata),  //       .writedata
		.byteenable (mm_interconnect_0_onchip_memory_s1_byteenable), //       .byteenable
		.reset      (rst_controller_001_reset_out_reset),            // reset1.reset
		.reset_req  (rst_controller_001_reset_out_reset_req),        //       .reset_req
		.freeze     (1'b0)                                           // (terminated)
	);

	NIOS_LED_Qsys_pll pll (
		.refclk   (clk_clk),         //  refclk.clk
		.rst      (~reset_reset_n),  //   reset.reset
		.outclk_0 (pll_outclk0_clk), // outclk0.clk
		.outclk_1 (pll_outclk1_clk), // outclk1.clk
		.locked   ()                 // (terminated)
	);

	NIOS_LED_Qsys_sysid sysid (
		.clock    (pll_outclk1_clk),                                //           clk.clk
		.reset_n  (~rst_controller_002_reset_out_reset),            //         reset.reset_n
		.readdata (mm_interconnect_1_sysid_control_slave_readdata), // control_slave.readdata
		.address  (mm_interconnect_1_sysid_control_slave_address)   //              .address
	);

	NIOS_LED_Qsys_timer_10ms timer_10ms (
		.clk        (pll_outclk1_clk),                            //   clk.clk
		.reset_n    (~rst_controller_002_reset_out_reset),        // reset.reset_n
		.address    (mm_interconnect_1_timer_10ms_s1_address),    //    s1.address
		.writedata  (mm_interconnect_1_timer_10ms_s1_writedata),  //      .writedata
		.readdata   (mm_interconnect_1_timer_10ms_s1_readdata),   //      .readdata
		.chipselect (mm_interconnect_1_timer_10ms_s1_chipselect), //      .chipselect
		.write_n    (~mm_interconnect_1_timer_10ms_s1_write),     //      .write_n
		.irq        (irq_synchronizer_001_receiver_irq)           //   irq.irq
	);

	NIOS_LED_Qsys_timer_1ms timer_1ms (
		.clk        (pll_outclk1_clk),                           //   clk.clk
		.reset_n    (~rst_controller_002_reset_out_reset),       // reset.reset_n
		.address    (mm_interconnect_1_timer_1ms_s1_address),    //    s1.address
		.writedata  (mm_interconnect_1_timer_1ms_s1_writedata),  //      .writedata
		.readdata   (mm_interconnect_1_timer_1ms_s1_readdata),   //      .readdata
		.chipselect (mm_interconnect_1_timer_1ms_s1_chipselect), //      .chipselect
		.write_n    (~mm_interconnect_1_timer_1ms_s1_write),     //      .write_n
		.irq        (irq_synchronizer_receiver_irq)              //   irq.irq
	);

	NIOS_LED_Qsys_mm_interconnect_0 mm_interconnect_0 (
		.pll_outclk0_clk                                               (pll_outclk0_clk),                                             //                                             pll_outclk0.clk
		.pll_outclk1_clk                                               (pll_outclk1_clk),                                             //                                             pll_outclk1.clk
		.mm_clock_crossing_bridge_s0_reset_reset_bridge_in_reset_reset (rst_controller_002_reset_out_reset),                          // mm_clock_crossing_bridge_s0_reset_reset_bridge_in_reset.reset
		.NIOS_CPU_reset_reset_bridge_in_reset_reset                    (rst_controller_001_reset_out_reset),                          //                    NIOS_CPU_reset_reset_bridge_in_reset.reset
		.NIOS_CPU_data_master_address                                  (nios_cpu_data_master_address),                                //                                    NIOS_CPU_data_master.address
		.NIOS_CPU_data_master_waitrequest                              (nios_cpu_data_master_waitrequest),                            //                                                        .waitrequest
		.NIOS_CPU_data_master_byteenable                               (nios_cpu_data_master_byteenable),                             //                                                        .byteenable
		.NIOS_CPU_data_master_read                                     (nios_cpu_data_master_read),                                   //                                                        .read
		.NIOS_CPU_data_master_readdata                                 (nios_cpu_data_master_readdata),                               //                                                        .readdata
		.NIOS_CPU_data_master_write                                    (nios_cpu_data_master_write),                                  //                                                        .write
		.NIOS_CPU_data_master_writedata                                (nios_cpu_data_master_writedata),                              //                                                        .writedata
		.NIOS_CPU_data_master_debugaccess                              (nios_cpu_data_master_debugaccess),                            //                                                        .debugaccess
		.NIOS_CPU_instruction_master_address                           (nios_cpu_instruction_master_address),                         //                             NIOS_CPU_instruction_master.address
		.NIOS_CPU_instruction_master_waitrequest                       (nios_cpu_instruction_master_waitrequest),                     //                                                        .waitrequest
		.NIOS_CPU_instruction_master_read                              (nios_cpu_instruction_master_read),                            //                                                        .read
		.NIOS_CPU_instruction_master_readdata                          (nios_cpu_instruction_master_readdata),                        //                                                        .readdata
		.mm_clock_crossing_bridge_s0_address                           (mm_interconnect_0_mm_clock_crossing_bridge_s0_address),       //                             mm_clock_crossing_bridge_s0.address
		.mm_clock_crossing_bridge_s0_write                             (mm_interconnect_0_mm_clock_crossing_bridge_s0_write),         //                                                        .write
		.mm_clock_crossing_bridge_s0_read                              (mm_interconnect_0_mm_clock_crossing_bridge_s0_read),          //                                                        .read
		.mm_clock_crossing_bridge_s0_readdata                          (mm_interconnect_0_mm_clock_crossing_bridge_s0_readdata),      //                                                        .readdata
		.mm_clock_crossing_bridge_s0_writedata                         (mm_interconnect_0_mm_clock_crossing_bridge_s0_writedata),     //                                                        .writedata
		.mm_clock_crossing_bridge_s0_burstcount                        (mm_interconnect_0_mm_clock_crossing_bridge_s0_burstcount),    //                                                        .burstcount
		.mm_clock_crossing_bridge_s0_byteenable                        (mm_interconnect_0_mm_clock_crossing_bridge_s0_byteenable),    //                                                        .byteenable
		.mm_clock_crossing_bridge_s0_readdatavalid                     (mm_interconnect_0_mm_clock_crossing_bridge_s0_readdatavalid), //                                                        .readdatavalid
		.mm_clock_crossing_bridge_s0_waitrequest                       (mm_interconnect_0_mm_clock_crossing_bridge_s0_waitrequest),   //                                                        .waitrequest
		.mm_clock_crossing_bridge_s0_debugaccess                       (mm_interconnect_0_mm_clock_crossing_bridge_s0_debugaccess),   //                                                        .debugaccess
		.NIOS_CPU_debug_mem_slave_address                              (mm_interconnect_0_nios_cpu_debug_mem_slave_address),          //                                NIOS_CPU_debug_mem_slave.address
		.NIOS_CPU_debug_mem_slave_write                                (mm_interconnect_0_nios_cpu_debug_mem_slave_write),            //                                                        .write
		.NIOS_CPU_debug_mem_slave_read                                 (mm_interconnect_0_nios_cpu_debug_mem_slave_read),             //                                                        .read
		.NIOS_CPU_debug_mem_slave_readdata                             (mm_interconnect_0_nios_cpu_debug_mem_slave_readdata),         //                                                        .readdata
		.NIOS_CPU_debug_mem_slave_writedata                            (mm_interconnect_0_nios_cpu_debug_mem_slave_writedata),        //                                                        .writedata
		.NIOS_CPU_debug_mem_slave_byteenable                           (mm_interconnect_0_nios_cpu_debug_mem_slave_byteenable),       //                                                        .byteenable
		.NIOS_CPU_debug_mem_slave_waitrequest                          (mm_interconnect_0_nios_cpu_debug_mem_slave_waitrequest),      //                                                        .waitrequest
		.NIOS_CPU_debug_mem_slave_debugaccess                          (mm_interconnect_0_nios_cpu_debug_mem_slave_debugaccess),      //                                                        .debugaccess
		.onchip_memory_s1_address                                      (mm_interconnect_0_onchip_memory_s1_address),                  //                                        onchip_memory_s1.address
		.onchip_memory_s1_write                                        (mm_interconnect_0_onchip_memory_s1_write),                    //                                                        .write
		.onchip_memory_s1_readdata                                     (mm_interconnect_0_onchip_memory_s1_readdata),                 //                                                        .readdata
		.onchip_memory_s1_writedata                                    (mm_interconnect_0_onchip_memory_s1_writedata),                //                                                        .writedata
		.onchip_memory_s1_byteenable                                   (mm_interconnect_0_onchip_memory_s1_byteenable),               //                                                        .byteenable
		.onchip_memory_s1_chipselect                                   (mm_interconnect_0_onchip_memory_s1_chipselect),               //                                                        .chipselect
		.onchip_memory_s1_clken                                        (mm_interconnect_0_onchip_memory_s1_clken)                     //                                                        .clken
	);

	NIOS_LED_Qsys_mm_interconnect_1 mm_interconnect_1 (
		.pll_outclk0_clk                                               (pll_outclk0_clk),                                           //                                             pll_outclk0.clk
		.pll_outclk1_clk                                               (pll_outclk1_clk),                                           //                                             pll_outclk1.clk
		.jtag_uart_reset_reset_bridge_in_reset_reset                   (rst_controller_001_reset_out_reset),                        //                   jtag_uart_reset_reset_bridge_in_reset.reset
		.LED_reset_reset_bridge_in_reset_reset                         (rst_controller_reset_out_reset),                            //                         LED_reset_reset_bridge_in_reset.reset
		.mm_clock_crossing_bridge_m0_reset_reset_bridge_in_reset_reset (rst_controller_002_reset_out_reset),                        // mm_clock_crossing_bridge_m0_reset_reset_bridge_in_reset.reset
		.mm_clock_crossing_bridge_m0_address                           (mm_clock_crossing_bridge_m0_address),                       //                             mm_clock_crossing_bridge_m0.address
		.mm_clock_crossing_bridge_m0_waitrequest                       (mm_clock_crossing_bridge_m0_waitrequest),                   //                                                        .waitrequest
		.mm_clock_crossing_bridge_m0_burstcount                        (mm_clock_crossing_bridge_m0_burstcount),                    //                                                        .burstcount
		.mm_clock_crossing_bridge_m0_byteenable                        (mm_clock_crossing_bridge_m0_byteenable),                    //                                                        .byteenable
		.mm_clock_crossing_bridge_m0_read                              (mm_clock_crossing_bridge_m0_read),                          //                                                        .read
		.mm_clock_crossing_bridge_m0_readdata                          (mm_clock_crossing_bridge_m0_readdata),                      //                                                        .readdata
		.mm_clock_crossing_bridge_m0_readdatavalid                     (mm_clock_crossing_bridge_m0_readdatavalid),                 //                                                        .readdatavalid
		.mm_clock_crossing_bridge_m0_write                             (mm_clock_crossing_bridge_m0_write),                         //                                                        .write
		.mm_clock_crossing_bridge_m0_writedata                         (mm_clock_crossing_bridge_m0_writedata),                     //                                                        .writedata
		.mm_clock_crossing_bridge_m0_debugaccess                       (mm_clock_crossing_bridge_m0_debugaccess),                   //                                                        .debugaccess
		.jtag_uart_avalon_jtag_slave_address                           (mm_interconnect_1_jtag_uart_avalon_jtag_slave_address),     //                             jtag_uart_avalon_jtag_slave.address
		.jtag_uart_avalon_jtag_slave_write                             (mm_interconnect_1_jtag_uart_avalon_jtag_slave_write),       //                                                        .write
		.jtag_uart_avalon_jtag_slave_read                              (mm_interconnect_1_jtag_uart_avalon_jtag_slave_read),        //                                                        .read
		.jtag_uart_avalon_jtag_slave_readdata                          (mm_interconnect_1_jtag_uart_avalon_jtag_slave_readdata),    //                                                        .readdata
		.jtag_uart_avalon_jtag_slave_writedata                         (mm_interconnect_1_jtag_uart_avalon_jtag_slave_writedata),   //                                                        .writedata
		.jtag_uart_avalon_jtag_slave_waitrequest                       (mm_interconnect_1_jtag_uart_avalon_jtag_slave_waitrequest), //                                                        .waitrequest
		.jtag_uart_avalon_jtag_slave_chipselect                        (mm_interconnect_1_jtag_uart_avalon_jtag_slave_chipselect),  //                                                        .chipselect
		.LED_s1_address                                                (mm_interconnect_1_led_s1_address),                          //                                                  LED_s1.address
		.LED_s1_write                                                  (mm_interconnect_1_led_s1_write),                            //                                                        .write
		.LED_s1_readdata                                               (mm_interconnect_1_led_s1_readdata),                         //                                                        .readdata
		.LED_s1_writedata                                              (mm_interconnect_1_led_s1_writedata),                        //                                                        .writedata
		.LED_s1_chipselect                                             (mm_interconnect_1_led_s1_chipselect),                       //                                                        .chipselect
		.SW_s1_address                                                 (mm_interconnect_1_sw_s1_address),                           //                                                   SW_s1.address
		.SW_s1_readdata                                                (mm_interconnect_1_sw_s1_readdata),                          //                                                        .readdata
		.sysid_control_slave_address                                   (mm_interconnect_1_sysid_control_slave_address),             //                                     sysid_control_slave.address
		.sysid_control_slave_readdata                                  (mm_interconnect_1_sysid_control_slave_readdata),            //                                                        .readdata
		.timer_10ms_s1_address                                         (mm_interconnect_1_timer_10ms_s1_address),                   //                                           timer_10ms_s1.address
		.timer_10ms_s1_write                                           (mm_interconnect_1_timer_10ms_s1_write),                     //                                                        .write
		.timer_10ms_s1_readdata                                        (mm_interconnect_1_timer_10ms_s1_readdata),                  //                                                        .readdata
		.timer_10ms_s1_writedata                                       (mm_interconnect_1_timer_10ms_s1_writedata),                 //                                                        .writedata
		.timer_10ms_s1_chipselect                                      (mm_interconnect_1_timer_10ms_s1_chipselect),                //                                                        .chipselect
		.timer_1ms_s1_address                                          (mm_interconnect_1_timer_1ms_s1_address),                    //                                            timer_1ms_s1.address
		.timer_1ms_s1_write                                            (mm_interconnect_1_timer_1ms_s1_write),                      //                                                        .write
		.timer_1ms_s1_readdata                                         (mm_interconnect_1_timer_1ms_s1_readdata),                   //                                                        .readdata
		.timer_1ms_s1_writedata                                        (mm_interconnect_1_timer_1ms_s1_writedata),                  //                                                        .writedata
		.timer_1ms_s1_chipselect                                       (mm_interconnect_1_timer_1ms_s1_chipselect)                  //                                                        .chipselect
	);

	NIOS_LED_Qsys_irq_mapper irq_mapper (
		.clk           (pll_outclk0_clk),                    //       clk.clk
		.reset         (rst_controller_001_reset_out_reset), // clk_reset.reset
		.receiver0_irq (irq_mapper_receiver0_irq),           // receiver0.irq
		.receiver1_irq (irq_mapper_receiver1_irq),           // receiver1.irq
		.receiver2_irq (irq_mapper_receiver2_irq),           // receiver2.irq
		.sender_irq    (nios_cpu_irq_irq)                    //    sender.irq
	);

	altera_irq_clock_crosser #(
		.IRQ_WIDTH (1)
	) irq_synchronizer (
		.receiver_clk   (pll_outclk1_clk),                    //       receiver_clk.clk
		.sender_clk     (pll_outclk0_clk),                    //         sender_clk.clk
		.receiver_reset (rst_controller_002_reset_out_reset), // receiver_clk_reset.reset
		.sender_reset   (rst_controller_001_reset_out_reset), //   sender_clk_reset.reset
		.receiver_irq   (irq_synchronizer_receiver_irq),      //           receiver.irq
		.sender_irq     (irq_mapper_receiver0_irq)            //             sender.irq
	);

	altera_irq_clock_crosser #(
		.IRQ_WIDTH (1)
	) irq_synchronizer_001 (
		.receiver_clk   (pll_outclk1_clk),                    //       receiver_clk.clk
		.sender_clk     (pll_outclk0_clk),                    //         sender_clk.clk
		.receiver_reset (rst_controller_002_reset_out_reset), // receiver_clk_reset.reset
		.sender_reset   (rst_controller_001_reset_out_reset), //   sender_clk_reset.reset
		.receiver_irq   (irq_synchronizer_001_receiver_irq),  //           receiver.irq
		.sender_irq     (irq_mapper_receiver1_irq)            //             sender.irq
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (1),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (0),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller (
		.reset_in0      (nios_cpu_debug_reset_request_reset), // reset_in0.reset
		.clk            (pll_outclk1_clk),                    //       clk.clk
		.reset_out      (rst_controller_reset_out_reset),     // reset_out.reset
		.reset_req      (),                                   // (terminated)
		.reset_req_in0  (1'b0),                               // (terminated)
		.reset_in1      (1'b0),                               // (terminated)
		.reset_req_in1  (1'b0),                               // (terminated)
		.reset_in2      (1'b0),                               // (terminated)
		.reset_req_in2  (1'b0),                               // (terminated)
		.reset_in3      (1'b0),                               // (terminated)
		.reset_req_in3  (1'b0),                               // (terminated)
		.reset_in4      (1'b0),                               // (terminated)
		.reset_req_in4  (1'b0),                               // (terminated)
		.reset_in5      (1'b0),                               // (terminated)
		.reset_req_in5  (1'b0),                               // (terminated)
		.reset_in6      (1'b0),                               // (terminated)
		.reset_req_in6  (1'b0),                               // (terminated)
		.reset_in7      (1'b0),                               // (terminated)
		.reset_req_in7  (1'b0),                               // (terminated)
		.reset_in8      (1'b0),                               // (terminated)
		.reset_req_in8  (1'b0),                               // (terminated)
		.reset_in9      (1'b0),                               // (terminated)
		.reset_req_in9  (1'b0),                               // (terminated)
		.reset_in10     (1'b0),                               // (terminated)
		.reset_req_in10 (1'b0),                               // (terminated)
		.reset_in11     (1'b0),                               // (terminated)
		.reset_req_in11 (1'b0),                               // (terminated)
		.reset_in12     (1'b0),                               // (terminated)
		.reset_req_in12 (1'b0),                               // (terminated)
		.reset_in13     (1'b0),                               // (terminated)
		.reset_req_in13 (1'b0),                               // (terminated)
		.reset_in14     (1'b0),                               // (terminated)
		.reset_req_in14 (1'b0),                               // (terminated)
		.reset_in15     (1'b0),                               // (terminated)
		.reset_req_in15 (1'b0)                                // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (2),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (1),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller_001 (
		.reset_in0      (~reset_reset_n),                         // reset_in0.reset
		.reset_in1      (nios_cpu_debug_reset_request_reset),     // reset_in1.reset
		.clk            (pll_outclk0_clk),                        //       clk.clk
		.reset_out      (rst_controller_001_reset_out_reset),     // reset_out.reset
		.reset_req      (rst_controller_001_reset_out_reset_req), //          .reset_req
		.reset_req_in0  (1'b0),                                   // (terminated)
		.reset_req_in1  (1'b0),                                   // (terminated)
		.reset_in2      (1'b0),                                   // (terminated)
		.reset_req_in2  (1'b0),                                   // (terminated)
		.reset_in3      (1'b0),                                   // (terminated)
		.reset_req_in3  (1'b0),                                   // (terminated)
		.reset_in4      (1'b0),                                   // (terminated)
		.reset_req_in4  (1'b0),                                   // (terminated)
		.reset_in5      (1'b0),                                   // (terminated)
		.reset_req_in5  (1'b0),                                   // (terminated)
		.reset_in6      (1'b0),                                   // (terminated)
		.reset_req_in6  (1'b0),                                   // (terminated)
		.reset_in7      (1'b0),                                   // (terminated)
		.reset_req_in7  (1'b0),                                   // (terminated)
		.reset_in8      (1'b0),                                   // (terminated)
		.reset_req_in8  (1'b0),                                   // (terminated)
		.reset_in9      (1'b0),                                   // (terminated)
		.reset_req_in9  (1'b0),                                   // (terminated)
		.reset_in10     (1'b0),                                   // (terminated)
		.reset_req_in10 (1'b0),                                   // (terminated)
		.reset_in11     (1'b0),                                   // (terminated)
		.reset_req_in11 (1'b0),                                   // (terminated)
		.reset_in12     (1'b0),                                   // (terminated)
		.reset_req_in12 (1'b0),                                   // (terminated)
		.reset_in13     (1'b0),                                   // (terminated)
		.reset_req_in13 (1'b0),                                   // (terminated)
		.reset_in14     (1'b0),                                   // (terminated)
		.reset_req_in14 (1'b0),                                   // (terminated)
		.reset_in15     (1'b0),                                   // (terminated)
		.reset_req_in15 (1'b0)                                    // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (2),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (0),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller_002 (
		.reset_in0      (~reset_reset_n),                     // reset_in0.reset
		.reset_in1      (nios_cpu_debug_reset_request_reset), // reset_in1.reset
		.clk            (pll_outclk1_clk),                    //       clk.clk
		.reset_out      (rst_controller_002_reset_out_reset), // reset_out.reset
		.reset_req      (),                                   // (terminated)
		.reset_req_in0  (1'b0),                               // (terminated)
		.reset_req_in1  (1'b0),                               // (terminated)
		.reset_in2      (1'b0),                               // (terminated)
		.reset_req_in2  (1'b0),                               // (terminated)
		.reset_in3      (1'b0),                               // (terminated)
		.reset_req_in3  (1'b0),                               // (terminated)
		.reset_in4      (1'b0),                               // (terminated)
		.reset_req_in4  (1'b0),                               // (terminated)
		.reset_in5      (1'b0),                               // (terminated)
		.reset_req_in5  (1'b0),                               // (terminated)
		.reset_in6      (1'b0),                               // (terminated)
		.reset_req_in6  (1'b0),                               // (terminated)
		.reset_in7      (1'b0),                               // (terminated)
		.reset_req_in7  (1'b0),                               // (terminated)
		.reset_in8      (1'b0),                               // (terminated)
		.reset_req_in8  (1'b0),                               // (terminated)
		.reset_in9      (1'b0),                               // (terminated)
		.reset_req_in9  (1'b0),                               // (terminated)
		.reset_in10     (1'b0),                               // (terminated)
		.reset_req_in10 (1'b0),                               // (terminated)
		.reset_in11     (1'b0),                               // (terminated)
		.reset_req_in11 (1'b0),                               // (terminated)
		.reset_in12     (1'b0),                               // (terminated)
		.reset_req_in12 (1'b0),                               // (terminated)
		.reset_in13     (1'b0),                               // (terminated)
		.reset_req_in13 (1'b0),                               // (terminated)
		.reset_in14     (1'b0),                               // (terminated)
		.reset_req_in14 (1'b0),                               // (terminated)
		.reset_in15     (1'b0),                               // (terminated)
		.reset_req_in15 (1'b0)                                // (terminated)
	);

endmodule
